library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;


entity WS2812_LED is
port (
	clk : in std_logic;
	reset : in std_logic;
	dout : out std_logic
	);
end WS2812_LED;

architecture behavior of WS2812_LED is

begin
	
		

end behavior;
